// decoder for nes controller