//My top level module for signal generation. Not much to see here honestly.
module signalgenerator(	input logic [8:0] keys,
						input logic reset,
						output logic [7:0] signal);
		
		logic clk;
		logic LUTclk;
		logic LUTsignal;
		
	//This is one of those magical built in modules that SystemVerilog gives us	
	OSCH #("2.08") osc_int (	//"2.08" specifies the operating frequency, 2.08 MHz.
									//Other clock frequencies can be found in the MachX02's documentation
			.STDBY(1'b0),			//Specifies active state
			.OSC(clk),				//Outputs clock signal to 'clk' net
			.SEDSTDBY());			//Leaves SEDSTDBY pin unconnected
	
	SignalClockDivider(	
			.keys(keys),
			.clk(clk),
			.signalLUTclk(LUTclk));
			
	SignalLUT(	
			.clk(LUTclk),
			.reset(reset),
			.signal(LUTsignal));
	
endmodule