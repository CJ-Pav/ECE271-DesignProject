// decoder for nes controller

