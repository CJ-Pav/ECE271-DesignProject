module signalLUT(	input logic clk, reset,
					output logic [7:0] signal
					);
	int counter;
	always_ff @(posedge clk, posedge reset)
			if (reset) counter <= 0;
			else if (counter == 524) counter <= 0;
			else counter <= counter + 1; 
	always_comb
		case(counter)
			0: signal <= 8'b10000000;
			1: signal <= 8'b10000001;
			2: signal <= 8'b10000011;
			3: signal <= 8'b10000100;
			4: signal <= 8'b10000110;
			5: signal <= 8'b10000111;
			6: signal <= 8'b10001001;
			7: signal <= 8'b10001010;
			8: signal <= 8'b10001100;
			9: signal <= 8'b10001101;
			10: signal <= 8'b10001111;
			11: signal <= 8'b10010000;
			12: signal <= 8'b10010010;
			13: signal <= 8'b10010011;
			14: signal <= 8'b10010101;
			15: signal <= 8'b10010110;
			16: signal <= 8'b10011000;
			17: signal <= 8'b10011001;
			18: signal <= 8'b10011011;
			19: signal <= 8'b10011100;
			20: signal <= 8'b10011110;
			21: signal <= 8'b10011111;
			22: signal <= 8'b10100001;
			23: signal <= 8'b10100010;
			24: signal <= 8'b10100100;
			25: signal <= 8'b10100101;
			26: signal <= 8'b10100111;
			27: signal <= 8'b10101000;
			28: signal <= 8'b10101010;
			29: signal <= 8'b10101011;
			30: signal <= 8'b10101100;
			31: signal <= 8'b10101110;
			32: signal <= 8'b10101111;
			33: signal <= 8'b10110001;
			34: signal <= 8'b10110010;
			35: signal <= 8'b10110100;
			36: signal <= 8'b10110101;
			37: signal <= 8'b10110110;
			38: signal <= 8'b10111000;
			39: signal <= 8'b10111001;
			40: signal <= 8'b10111010;
			41: signal <= 8'b10111100;
			42: signal <= 8'b10111101;
			43: signal <= 8'b10111111;
			44: signal <= 8'b11000000;
			45: signal <= 8'b11000001;
			46: signal <= 8'b11000010;
			47: signal <= 8'b11000100;
			48: signal <= 8'b11000101;
			49: signal <= 8'b11000110;
			50: signal <= 8'b11001000;
			51: signal <= 8'b11001001;
			52: signal <= 8'b11001010;
			53: signal <= 8'b11001011;
			54: signal <= 8'b11001101;
			55: signal <= 8'b11001110;
			56: signal <= 8'b11001111;
			57: signal <= 8'b11010000;
			58: signal <= 8'b11010001;
			59: signal <= 8'b11010011;
			60: signal <= 8'b11010100;
			61: signal <= 8'b11010101;
			62: signal <= 8'b11010110;
			63: signal <= 8'b11010111;
			64: signal <= 8'b11011000;
			65: signal <= 8'b11011001;
			66: signal <= 8'b11011010;
			67: signal <= 8'b11011011;
			68: signal <= 8'b11011101;
			69: signal <= 8'b11011110;
			70: signal <= 8'b11011111;
			71: signal <= 8'b11100000;
			72: signal <= 8'b11100001;
			73: signal <= 8'b11100010;
			74: signal <= 8'b11100011;
			75: signal <= 8'b11100100;
			76: signal <= 8'b11100101;
			77: signal <= 8'b11100101;
			78: signal <= 8'b11100110;
			79: signal <= 8'b11100111;
			80: signal <= 8'b11101000;
			81: signal <= 8'b11101001;
			82: signal <= 8'b11101010;
			83: signal <= 8'b11101011;
			84: signal <= 8'b11101100;
			85: signal <= 8'b11101100;
			86: signal <= 8'b11101101;
			87: signal <= 8'b11101110;
			88: signal <= 8'b11101111;
			89: signal <= 8'b11101111;
			90: signal <= 8'b11110000;
			91: signal <= 8'b11110001;
			92: signal <= 8'b11110010;
			93: signal <= 8'b11110010;
			94: signal <= 8'b11110011;
			95: signal <= 8'b11110100;
			96: signal <= 8'b11110100;
			97: signal <= 8'b11110101;
			98: signal <= 8'b11110101;
			99: signal <= 8'b11110110;
			100: signal <= 8'b11110111;
			101: signal <= 8'b11110111;
			102: signal <= 8'b11111000;
			103: signal <= 8'b11111000;
			104: signal <= 8'b11111001;
			105: signal <= 8'b11111001;
			106: signal <= 8'b11111010;
			107: signal <= 8'b11111010;
			108: signal <= 8'b11111011;
			109: signal <= 8'b11111011;
			110: signal <= 8'b11111011;
			111: signal <= 8'b11111100;
			112: signal <= 8'b11111100;
			113: signal <= 8'b11111100;
			114: signal <= 8'b11111101;
			115: signal <= 8'b11111101;
			116: signal <= 8'b11111101;
			117: signal <= 8'b11111110;
			118: signal <= 8'b11111110;
			119: signal <= 8'b11111110;
			120: signal <= 8'b11111110;
			121: signal <= 8'b11111111;
			122: signal <= 8'b11111111;
			123: signal <= 8'b11111111;
			124: signal <= 8'b11111111;
			125: signal <= 8'b11111111;
			126: signal <= 8'b11111111;
			127: signal <= 8'b11111111;
			128: signal <= 8'b11111111;
			129: signal <= 8'b11111111;
			130: signal <= 8'b11111111;
			131: signal <= 8'b11111111;
			132: signal <= 8'b11111111;
			133: signal <= 8'b11111111;
			134: signal <= 8'b11111111;
			135: signal <= 8'b11111111;
			136: signal <= 8'b11111111;
			137: signal <= 8'b11111111;
			138: signal <= 8'b11111111;
			139: signal <= 8'b11111111;
			140: signal <= 8'b11111111;
			141: signal <= 8'b11111111;
			142: signal <= 8'b11111110;
			143: signal <= 8'b11111110;
			144: signal <= 8'b11111110;
			145: signal <= 8'b11111110;
			146: signal <= 8'b11111110;
			147: signal <= 8'b11111101;
			148: signal <= 8'b11111101;
			149: signal <= 8'b11111101;
			150: signal <= 8'b11111100;
			151: signal <= 8'b11111100;
			152: signal <= 8'b11111100;
			153: signal <= 8'b11111011;
			154: signal <= 8'b11111011;
			155: signal <= 8'b11111010;
			156: signal <= 8'b11111010;
			157: signal <= 8'b11111001;
			158: signal <= 8'b11111001;
			159: signal <= 8'b11111001;
			160: signal <= 8'b11111000;
			161: signal <= 8'b11110111;
			162: signal <= 8'b11110111;
			163: signal <= 8'b11110110;
			164: signal <= 8'b11110110;
			165: signal <= 8'b11110101;
			166: signal <= 8'b11110101;
			167: signal <= 8'b11110100;
			168: signal <= 8'b11110011;
			169: signal <= 8'b11110011;
			170: signal <= 8'b11110010;
			171: signal <= 8'b11110001;
			172: signal <= 8'b11110001;
			173: signal <= 8'b11110000;
			174: signal <= 8'b11101111;
			175: signal <= 8'b11101110;
			176: signal <= 8'b11101110;
			177: signal <= 8'b11101101;
			178: signal <= 8'b11101100;
			179: signal <= 8'b11101011;
			180: signal <= 8'b11101010;
			181: signal <= 8'b11101001;
			182: signal <= 8'b11101001;
			183: signal <= 8'b11101000;
			184: signal <= 8'b11100111;
			185: signal <= 8'b11100110;
			186: signal <= 8'b11100101;
			187: signal <= 8'b11100100;
			188: signal <= 8'b11100011;
			189: signal <= 8'b11100010;
			190: signal <= 8'b11100001;
			191: signal <= 8'b11100000;
			192: signal <= 8'b11011111;
			193: signal <= 8'b11011110;
			194: signal <= 8'b11011101;
			195: signal <= 8'b11011100;
			196: signal <= 8'b11011011;
			197: signal <= 8'b11011010;
			198: signal <= 8'b11011001;
			199: signal <= 8'b11011000;
			200: signal <= 8'b11010111;
			201: signal <= 8'b11010101;
			202: signal <= 8'b11010100;
			203: signal <= 8'b11010011;
			204: signal <= 8'b11010010;
			205: signal <= 8'b11010001;
			206: signal <= 8'b11010000;
			207: signal <= 8'b11001110;
			208: signal <= 8'b11001101;
			209: signal <= 8'b11001100;
			210: signal <= 8'b11001011;
			211: signal <= 8'b11001001;
			212: signal <= 8'b11001000;
			213: signal <= 8'b11000111;
			214: signal <= 8'b11000110;
			215: signal <= 8'b11000100;
			216: signal <= 8'b11000011;
			217: signal <= 8'b11000010;
			218: signal <= 8'b11000000;
			219: signal <= 8'b10111111;
			220: signal <= 8'b10111110;
			221: signal <= 8'b10111100;
			222: signal <= 8'b10111011;
			223: signal <= 8'b10111010;
			224: signal <= 8'b10111000;
			225: signal <= 8'b10110111;
			226: signal <= 8'b10110110;
			227: signal <= 8'b10110100;
			228: signal <= 8'b10110011;
			229: signal <= 8'b10110001;
			230: signal <= 8'b10110000;
			231: signal <= 8'b10101111;
			232: signal <= 8'b10101101;
			233: signal <= 8'b10101100;
			234: signal <= 8'b10101010;
			235: signal <= 8'b10101001;
			236: signal <= 8'b10100111;
			237: signal <= 8'b10100110;
			238: signal <= 8'b10100100;
			239: signal <= 8'b10100011;
			240: signal <= 8'b10100010;
			241: signal <= 8'b10100000;
			242: signal <= 8'b10011111;
			243: signal <= 8'b10011101;
			244: signal <= 8'b10011100;
			245: signal <= 8'b10011010;
			246: signal <= 8'b10011001;
			247: signal <= 8'b10010111;
			248: signal <= 8'b10010110;
			249: signal <= 8'b10010100;
			250: signal <= 8'b10010011;
			251: signal <= 8'b10010001;
			252: signal <= 8'b10010000;
			253: signal <= 8'b10001110;
			254: signal <= 8'b10001100;
			255: signal <= 8'b10001011;
			256: signal <= 8'b10001001;
			257: signal <= 8'b10001000;
			258: signal <= 8'b10000110;
			259: signal <= 8'b10000101;
			260: signal <= 8'b10000011;
			261: signal <= 8'b10000010;
			262: signal <= 8'b10000000;
			263: signal <= 8'b01111111;
			264: signal <= 8'b01111101;
			265: signal <= 8'b01111100;
			266: signal <= 8'b01111010;
			267: signal <= 8'b01111001;
			268: signal <= 8'b01110111;
			269: signal <= 8'b01110110;
			270: signal <= 8'b01110100;
			271: signal <= 8'b01110010;
			272: signal <= 8'b01110001;
			273: signal <= 8'b01101111;
			274: signal <= 8'b01101110;
			275: signal <= 8'b01101100;
			276: signal <= 8'b01101011;
			277: signal <= 8'b01101001;
			278: signal <= 8'b01101000;
			279: signal <= 8'b01100110;
			280: signal <= 8'b01100101;
			281: signal <= 8'b01100011;
			282: signal <= 8'b01100010;
			283: signal <= 8'b01100000;
			284: signal <= 8'b01011111;
			285: signal <= 8'b01011101;
			286: signal <= 8'b01011100;
			287: signal <= 8'b01011011;
			288: signal <= 8'b01011001;
			289: signal <= 8'b01011000;
			290: signal <= 8'b01010110;
			291: signal <= 8'b01010101;
			292: signal <= 8'b01010011;
			293: signal <= 8'b01010010;
			294: signal <= 8'b01010000;
			295: signal <= 8'b01001111;
			296: signal <= 8'b01001110;
			297: signal <= 8'b01001100;
			298: signal <= 8'b01001011;
			299: signal <= 8'b01001001;
			300: signal <= 8'b01001000;
			301: signal <= 8'b01000111;
			302: signal <= 8'b01000101;
			303: signal <= 8'b01000100;
			304: signal <= 8'b01000011;
			305: signal <= 8'b01000001;
			306: signal <= 8'b01000000;
			307: signal <= 8'b00111111;
			308: signal <= 8'b00111101;
			309: signal <= 8'b00111100;
			310: signal <= 8'b00111011;
			311: signal <= 8'b00111001;
			312: signal <= 8'b00111000;
			313: signal <= 8'b00110111;
			314: signal <= 8'b00110110;
			315: signal <= 8'b00110100;
			316: signal <= 8'b00110011;
			317: signal <= 8'b00110010;
			318: signal <= 8'b00110001;
			319: signal <= 8'b00101111;
			320: signal <= 8'b00101110;
			321: signal <= 8'b00101101;
			322: signal <= 8'b00101100;
			323: signal <= 8'b00101011;
			324: signal <= 8'b00101010;
			325: signal <= 8'b00101000;
			326: signal <= 8'b00100111;
			327: signal <= 8'b00100110;
			328: signal <= 8'b00100101;
			329: signal <= 8'b00100100;
			330: signal <= 8'b00100011;
			331: signal <= 8'b00100010;
			332: signal <= 8'b00100001;
			333: signal <= 8'b00100000;
			334: signal <= 8'b00011111;
			335: signal <= 8'b00011110;
			336: signal <= 8'b00011101;
			337: signal <= 8'b00011100;
			338: signal <= 8'b00011011;
			339: signal <= 8'b00011010;
			340: signal <= 8'b00011001;
			341: signal <= 8'b00011000;
			342: signal <= 8'b00010111;
			343: signal <= 8'b00010110;
			344: signal <= 8'b00010110;
			345: signal <= 8'b00010101;
			346: signal <= 8'b00010100;
			347: signal <= 8'b00010011;
			348: signal <= 8'b00010010;
			349: signal <= 8'b00010001;
			350: signal <= 8'b00010001;
			351: signal <= 8'b00010000;
			352: signal <= 8'b00001111;
			353: signal <= 8'b00001110;
			354: signal <= 8'b00001110;
			355: signal <= 8'b00001101;
			356: signal <= 8'b00001100;
			357: signal <= 8'b00001100;
			358: signal <= 8'b00001011;
			359: signal <= 8'b00001010;
			360: signal <= 8'b00001010;
			361: signal <= 8'b00001001;
			362: signal <= 8'b00001001;
			363: signal <= 8'b00001000;
			364: signal <= 8'b00001000;
			365: signal <= 8'b00000111;
			366: signal <= 8'b00000110;
			367: signal <= 8'b00000110;
			368: signal <= 8'b00000110;
			369: signal <= 8'b00000101;
			370: signal <= 8'b00000101;
			371: signal <= 8'b00000100;
			372: signal <= 8'b00000100;
			373: signal <= 8'b00000011;
			374: signal <= 8'b00000011;
			375: signal <= 8'b00000011;
			376: signal <= 8'b00000010;
			377: signal <= 8'b00000010;
			378: signal <= 8'b00000010;
			379: signal <= 8'b00000001;
			380: signal <= 8'b00000001;
			381: signal <= 8'b00000001;
			382: signal <= 8'b00000001;
			383: signal <= 8'b00000001;
			384: signal <= 8'b00000000;
			385: signal <= 8'b00000000;
			386: signal <= 8'b00000000;
			387: signal <= 8'b00000000;
			388: signal <= 8'b00000000;
			389: signal <= 8'b00000000;
			390: signal <= 8'b00000000;
			391: signal <= 8'b00000000;
			392: signal <= 8'b00000000;
			393: signal <= 8'b00000000;
			394: signal <= 8'b00000000;
			395: signal <= 8'b00000000;
			396: signal <= 8'b00000000;
			397: signal <= 8'b00000000;
			398: signal <= 8'b00000000;
			399: signal <= 8'b00000000;
			400: signal <= 8'b00000000;
			401: signal <= 8'b00000000;
			402: signal <= 8'b00000000;
			403: signal <= 8'b00000000;
			404: signal <= 8'b00000000;
			405: signal <= 8'b00000001;
			406: signal <= 8'b00000001;
			407: signal <= 8'b00000001;
			408: signal <= 8'b00000001;
			409: signal <= 8'b00000010;
			410: signal <= 8'b00000010;
			411: signal <= 8'b00000010;
			412: signal <= 8'b00000011;
			413: signal <= 8'b00000011;
			414: signal <= 8'b00000011;
			415: signal <= 8'b00000100;
			416: signal <= 8'b00000100;
			417: signal <= 8'b00000100;
			418: signal <= 8'b00000101;
			419: signal <= 8'b00000101;
			420: signal <= 8'b00000110;
			421: signal <= 8'b00000110;
			422: signal <= 8'b00000111;
			423: signal <= 8'b00000111;
			424: signal <= 8'b00001000;
			425: signal <= 8'b00001000;
			426: signal <= 8'b00001001;
			427: signal <= 8'b00001010;
			428: signal <= 8'b00001010;
			429: signal <= 8'b00001011;
			430: signal <= 8'b00001011;
			431: signal <= 8'b00001100;
			432: signal <= 8'b00001101;
			433: signal <= 8'b00001101;
			434: signal <= 8'b00001110;
			435: signal <= 8'b00001111;
			436: signal <= 8'b00010000;
			437: signal <= 8'b00010000;
			438: signal <= 8'b00010001;
			439: signal <= 8'b00010010;
			440: signal <= 8'b00010011;
			441: signal <= 8'b00010011;
			442: signal <= 8'b00010100;
			443: signal <= 8'b00010101;
			444: signal <= 8'b00010110;
			445: signal <= 8'b00010111;
			446: signal <= 8'b00011000;
			447: signal <= 8'b00011001;
			448: signal <= 8'b00011010;
			449: signal <= 8'b00011010;
			450: signal <= 8'b00011011;
			451: signal <= 8'b00011100;
			452: signal <= 8'b00011101;
			453: signal <= 8'b00011110;
			454: signal <= 8'b00011111;
			455: signal <= 8'b00100000;
			456: signal <= 8'b00100001;
			457: signal <= 8'b00100010;
			458: signal <= 8'b00100100;
			459: signal <= 8'b00100101;
			460: signal <= 8'b00100110;
			461: signal <= 8'b00100111;
			462: signal <= 8'b00101000;
			463: signal <= 8'b00101001;
			464: signal <= 8'b00101010;
			465: signal <= 8'b00101011;
			466: signal <= 8'b00101100;
			467: signal <= 8'b00101110;
			468: signal <= 8'b00101111;
			469: signal <= 8'b00110000;
			470: signal <= 8'b00110001;
			471: signal <= 8'b00110010;
			472: signal <= 8'b00110100;
			473: signal <= 8'b00110101;
			474: signal <= 8'b00110110;
			475: signal <= 8'b00110111;
			476: signal <= 8'b00111001;
			477: signal <= 8'b00111010;
			478: signal <= 8'b00111011;
			479: signal <= 8'b00111101;
			480: signal <= 8'b00111110;
			481: signal <= 8'b00111111;
			482: signal <= 8'b01000001;
			483: signal <= 8'b01000010;
			484: signal <= 8'b01000011;
			485: signal <= 8'b01000101;
			486: signal <= 8'b01000110;
			487: signal <= 8'b01000111;
			488: signal <= 8'b01001001;
			489: signal <= 8'b01001010;
			490: signal <= 8'b01001011;
			491: signal <= 8'b01001101;
			492: signal <= 8'b01001110;
			493: signal <= 8'b01010000;
			494: signal <= 8'b01010001;
			495: signal <= 8'b01010011;
			496: signal <= 8'b01010100;
			497: signal <= 8'b01010101;
			498: signal <= 8'b01010111;
			499: signal <= 8'b01011000;
			500: signal <= 8'b01011010;
			501: signal <= 8'b01011011;
			502: signal <= 8'b01011101;
			503: signal <= 8'b01011110;
			504: signal <= 8'b01100000;
			505: signal <= 8'b01100001;
			506: signal <= 8'b01100011;
			507: signal <= 8'b01100100;
			508: signal <= 8'b01100110;
			509: signal <= 8'b01100111;
			510: signal <= 8'b01101001;
			511: signal <= 8'b01101010;
			512: signal <= 8'b01101100;
			513: signal <= 8'b01101101;
			514: signal <= 8'b01101111;
			515: signal <= 8'b01110000;
			516: signal <= 8'b01110010;
			517: signal <= 8'b01110011;
			518: signal <= 8'b01110101;
			519: signal <= 8'b01110110;
			520: signal <= 8'b01111000;
			521: signal <= 8'b01111001;
			522: signal <= 8'b01111011;
			523: signal <= 8'b01111100;
			524: signal <= 8'b01111110;
		endcase
endmodule