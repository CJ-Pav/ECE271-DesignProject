// one module to rule them all...