//This module doesn't currently work. The output logic named
//"signal" is a binary variable, and I am trying to assign
//it a real number value. It gets this number and just rounds
//it down to zero. Need to talk to the TAs to fix this
//problem.

//Also, I am assuming that the default timescale is 1ns
//(which it may not be). I couldn't get the 'timescale
//directive to work, so I'm just hoping it will 1ns
//by default.

module signalgenerator(	input logic [8:0] keys,
						output real signal);
		logic timestep = 440;
	always_comb
		case(keys)
			9'b100000000: timestep = 10**9 / (261.63*1024);
			9'b010000000: timestep = 10**9 / (293.67*1024);
			9'b001000000: timestep = 10**9 / (329.63*1024);
			9'b100100000: timestep = 10**9 / (349.23*1024);
			9'b100010000: timestep = 10**9 / (391.00*1024);
			9'b100001000: timestep = 10**9 / (440.00*1024);
			9'b100000100: timestep = 10**9 / (493.88*1024);
			9'b100000010: timestep = 10**9 / (523.25*1024);
			9'b100000001: timestep = 999999999;
		endcase
	
	always 
		begin 
			signal=0.5; #timestep;
			signal=0.503068; #timestep;
			signal=0.506136; #timestep;
			signal=0.509204; #timestep;
			signal=0.512271; #timestep;
			signal=0.515338; #timestep;
			signal=0.518404; #timestep;
			signal=0.52147; #timestep;
			signal=0.524535; #timestep;
			signal=0.527598; #timestep;
			signal=0.530661; #timestep;
			signal=0.533723; #timestep;
			signal=0.536783; #timestep;
			signal=0.539842; #timestep;
			signal=0.5429; #timestep;
			signal=0.545956; #timestep;
			signal=0.54901; #timestep;
			signal=0.552062; #timestep;
			signal=0.555113; #timestep;
			signal=0.558161; #timestep;
			signal=0.561207; #timestep;
			signal=0.564251; #timestep;
			signal=0.567292; #timestep;
			signal=0.570331; #timestep;
			signal=0.573367; #timestep;
			signal=0.576401; #timestep;
			signal=0.579431; #timestep;
			signal=0.582459; #timestep;
			signal=0.585483; #timestep;
			signal=0.588505; #timestep;
			signal=0.591523; #timestep;
			signal=0.594537; #timestep;
			signal=0.597548; #timestep;
			signal=0.600555; #timestep;
			signal=0.603559; #timestep;
			signal=0.606558; #timestep;
			signal=0.609554; #timestep;
			signal=0.612545; #timestep;
			signal=0.615532; #timestep;
			signal=0.618515; #timestep;
			signal=0.621493; #timestep;
			signal=0.624467; #timestep;
			signal=0.627436; #timestep;
			signal=0.630401; #timestep;
			signal=0.63336; #timestep;
			signal=0.636314; #timestep;
			signal=0.639264; #timestep;
			signal=0.642208; #timestep;
			signal=0.645146; #timestep;
			signal=0.64808; #timestep;
			signal=0.651007; #timestep;
			signal=0.653929; #timestep;
			signal=0.656845; #timestep;
			signal=0.659755; #timestep;
			signal=0.66266; #timestep;
			signal=0.665558; #timestep;
			signal=0.66845; #timestep;
			signal=0.671335; #timestep;
			signal=0.674214; #timestep;
			signal=0.677087; #timestep;
			signal=0.679952; #timestep;
			signal=0.682811; #timestep;
			signal=0.685664; #timestep;
			signal=0.688509; #timestep;
			signal=0.691347; #timestep;
			signal=0.694178; #timestep;
			signal=0.697001; #timestep;
			signal=0.699817; #timestep;
			signal=0.702626; #timestep;
			signal=0.705427; #timestep;
			signal=0.70822; #timestep;
			signal=0.711006; #timestep;
			signal=0.713783; #timestep;
			signal=0.716553; #timestep;
			signal=0.719314; #timestep;
			signal=0.722067; #timestep;
			signal=0.724812; #timestep;
			signal=0.727548; #timestep;
			signal=0.730275; #timestep;
			signal=0.732994; #timestep;
			signal=0.735705; #timestep;
			signal=0.738406; #timestep;
			signal=0.741098; #timestep;
			signal=0.743781; #timestep;
			signal=0.746456; #timestep;
			signal=0.74912; #timestep;
			signal=0.751776; #timestep;
			signal=0.754422; #timestep;
			signal=0.757058; #timestep;
			signal=0.759685; #timestep;
			signal=0.762302; #timestep;
			signal=0.764909; #timestep;
			signal=0.767506; #timestep;
			signal=0.770093; #timestep;
			signal=0.772669; #timestep;
			signal=0.775236; #timestep;
			signal=0.777792; #timestep;
			signal=0.780338; #timestep;
			signal=0.782873; #timestep;
			signal=0.785398; #timestep;
			signal=0.787911; #timestep;
			signal=0.790414; #timestep;
			signal=0.792906; #timestep;
			signal=0.795387; #timestep;
			signal=0.797857; #timestep;
			signal=0.800316; #timestep;
			signal=0.802763; #timestep;
			signal=0.805199; #timestep;
			signal=0.807623; #timestep;
			signal=0.810036; #timestep;
			signal=0.812437; #timestep;
			signal=0.814827; #timestep;
			signal=0.817204; #timestep;
			signal=0.81957; #timestep;
			signal=0.821923; #timestep;
			signal=0.824265; #timestep;
			signal=0.826594; #timestep;
			signal=0.828911; #timestep;
			signal=0.831216; #timestep;
			signal=0.833508; #timestep;
			signal=0.835787; #timestep;
			signal=0.838054; #timestep;
			signal=0.840308; #timestep;
			signal=0.84255; #timestep;
			signal=0.844778; #timestep;
			signal=0.846994; #timestep;
			signal=0.849196; #timestep;
			signal=0.851385; #timestep;
			signal=0.853561; #timestep;
			signal=0.855724; #timestep;
			signal=0.857873; #timestep;
			signal=0.860009; #timestep;
			signal=0.862132; #timestep;
			signal=0.86424; #timestep;
			signal=0.866335; #timestep;
			signal=0.868416; #timestep;
			signal=0.870484; #timestep;
			signal=0.872537; #timestep;
			signal=0.874576; #timestep;
			signal=0.876601; #timestep;
			signal=0.878612; #timestep;
			signal=0.880609; #timestep;
			signal=0.882592; #timestep;
			signal=0.88456; #timestep;
			signal=0.886513; #timestep;
			signal=0.888452; #timestep;
			signal=0.890377; #timestep;
			signal=0.892286; #timestep;
			signal=0.894181; #timestep;
			signal=0.896061; #timestep;
			signal=0.897926; #timestep;
			signal=0.899777; #timestep;
			signal=0.901612; #timestep;
			signal=0.903432; #timestep;
			signal=0.905237; #timestep;
			signal=0.907026; #timestep;
			signal=0.9088; #timestep;
			signal=0.910559; #timestep;
			signal=0.912302; #timestep;
			signal=0.91403; #timestep;
			signal=0.915743; #timestep;
			signal=0.917439; #timestep;
			signal=0.91912; #timestep;
			signal=0.920785; #timestep;
			signal=0.922434; #timestep;
			signal=0.924068; #timestep;
			signal=0.925685; #timestep;
			signal=0.927287; #timestep;
			signal=0.928872; #timestep;
			signal=0.930441; #timestep;
			signal=0.931994; #timestep;
			signal=0.933531; #timestep;
			signal=0.935051; #timestep;
			signal=0.936555; #timestep;
			signal=0.938042; #timestep;
			signal=0.939513; #timestep;
			signal=0.940968; #timestep;
			signal=0.942406; #timestep;
			signal=0.943827; #timestep;
			signal=0.945232; #timestep;
			signal=0.946619; #timestep;
			signal=0.94799; #timestep;
			signal=0.949344; #timestep;
			signal=0.950681; #timestep;
			signal=0.952002; #timestep;
			signal=0.953305; #timestep;
			signal=0.954591; #timestep;
			signal=0.95586; #timestep;
			signal=0.957112; #timestep;
			signal=0.958346; #timestep;
			signal=0.959563; #timestep;
			signal=0.960764; #timestep;
			signal=0.961946; #timestep;
			signal=0.963112; #timestep;
			signal=0.964259; #timestep;
			signal=0.96539; #timestep;
			signal=0.966503; #timestep;
			signal=0.967598; #timestep;
			signal=0.968676; #timestep;
			signal=0.969736; #timestep;
			signal=0.970778; #timestep;
			signal=0.971803; #timestep;
			signal=0.972809; #timestep;
			signal=0.973798; #timestep;
			signal=0.97477; #timestep;
			signal=0.975723; #timestep;
			signal=0.976658; #timestep;
			signal=0.977576; #timestep;
			signal=0.978475; #timestep;
			signal=0.979357; #timestep;
			signal=0.98022; #timestep;
			signal=0.981066; #timestep;
			signal=0.981893; #timestep;
			signal=0.982702; #timestep;
			signal=0.983493; #timestep;
			signal=0.984266; #timestep;
			signal=0.98502; #timestep;
			signal=0.985756; #timestep;
			signal=0.986474; #timestep;
			signal=0.987174; #timestep;
			signal=0.987855; #timestep;
			signal=0.988518; #timestep;
			signal=0.989163; #timestep;
			signal=0.989789; #timestep;
			signal=0.990396; #timestep;
			signal=0.990986; #timestep;
			signal=0.991556; #timestep;
			signal=0.992109; #timestep;
			signal=0.992642; #timestep;
			signal=0.993157; #timestep;
			signal=0.993654; #timestep;
			signal=0.994132; #timestep;
			signal=0.994591; #timestep;
			signal=0.995032; #timestep;
			signal=0.995454; #timestep;
			signal=0.995858; #timestep;
			signal=0.996242; #timestep;
			signal=0.996608; #timestep;
			signal=0.996956; #timestep;
			signal=0.997284; #timestep;
			signal=0.997594; #timestep;
			signal=0.997886; #timestep;
			signal=0.998158; #timestep;
			signal=0.998412; #timestep;
			signal=0.998647; #timestep;
			signal=0.998863; #timestep;
			signal=0.99906; #timestep;
			signal=0.999239; #timestep;
			signal=0.999399; #timestep;
			signal=0.99954; #timestep;
			signal=0.999662; #timestep;
			signal=0.999765; #timestep;
			signal=0.99985; #timestep;
			signal=0.999916; #timestep;
			signal=0.999963; #timestep;
			signal=0.999991; #timestep;
			signal=1; #timestep;
			signal=0.99999; #timestep;
			signal=0.999962; #timestep;
			signal=0.999915; #timestep;
			signal=0.999849; #timestep;
			signal=0.999764; #timestep;
			signal=0.99966; #timestep;
			signal=0.999538; #timestep;
			signal=0.999397; #timestep;
			signal=0.999237; #timestep;
			signal=0.999058; #timestep;
			signal=0.99886; #timestep;
			signal=0.998643; #timestep;
			signal=0.998408; #timestep;
			signal=0.998154; #timestep;
			signal=0.997882; #timestep;
			signal=0.99759; #timestep;
			signal=0.99728; #timestep;
			signal=0.996951; #timestep;
			signal=0.996603; #timestep;
			signal=0.996237; #timestep;
			signal=0.995852; #timestep;
			signal=0.995448; #timestep;
			signal=0.995026; #timestep;
			signal=0.994585; #timestep;
			signal=0.994125; #timestep;
			signal=0.993647; #timestep;
			signal=0.99315; #timestep;
			signal=0.992635; #timestep;
			signal=0.992101; #timestep;
			signal=0.991548; #timestep;
			signal=0.990977; #timestep;
			signal=0.990388; #timestep;
			signal=0.98978; #timestep;
			signal=0.989153; #timestep;
			signal=0.988509; #timestep;
			signal=0.987845; #timestep;
			signal=0.987164; #timestep;
			signal=0.986464; #timestep;
			signal=0.985746; #timestep;
			signal=0.985009; #timestep;
			signal=0.984255; #timestep;
			signal=0.983482; #timestep;
			signal=0.98269; #timestep;
			signal=0.981881; #timestep;
			signal=0.981054; #timestep;
			signal=0.980208; #timestep;
			signal=0.979344; #timestep;
			signal=0.978462; #timestep;
			signal=0.977563; #timestep;
			signal=0.976645; #timestep;
			signal=0.975709; #timestep;
			signal=0.974756; #timestep;
			signal=0.973784; #timestep;
			signal=0.972795; #timestep;
			signal=0.971788; #timestep;
			signal=0.970763; #timestep;
			signal=0.96972; #timestep;
			signal=0.96866; #timestep;
			signal=0.967582; #timestep;
			signal=0.966486; #timestep;
			signal=0.965373; #timestep;
			signal=0.964243; #timestep;
			signal=0.963095; #timestep;
			signal=0.961929; #timestep;
			signal=0.960746; #timestep;
			signal=0.959546; #timestep;
			signal=0.958328; #timestep;
			signal=0.957093; #timestep;
			signal=0.955841; #timestep;
			signal=0.954572; #timestep;
			signal=0.953286; #timestep;
			signal=0.951982; #timestep;
			signal=0.950662; #timestep;
			signal=0.949325; #timestep;
			signal=0.94797; #timestep;
			signal=0.946599; #timestep;
			signal=0.945211; #timestep;
			signal=0.943806; #timestep;
			signal=0.942385; #timestep;
			signal=0.940947; #timestep;
			signal=0.939492; #timestep;
			signal=0.938021; #timestep;
			signal=0.936533; #timestep;
			signal=0.935029; #timestep;
			signal=0.933508; #timestep;
			signal=0.931971; #timestep;
			signal=0.930418; #timestep;
			signal=0.928849; #timestep;
			signal=0.927263; #timestep;
			signal=0.925662; #timestep;
			signal=0.924044; #timestep;
			signal=0.92241; #timestep;
			signal=0.920761; #timestep;
			signal=0.919096; #timestep;
			signal=0.917414; #timestep;
			signal=0.915718; #timestep;
			signal=0.914005; #timestep;
			signal=0.912277; #timestep;
			signal=0.910533; #timestep;
			signal=0.908774; #timestep;
			signal=0.907; #timestep;
			signal=0.90521; #timestep;
			signal=0.903405; #timestep;
			signal=0.901585; #timestep;
			signal=0.89975; #timestep;
			signal=0.897899; #timestep;
			signal=0.896034; #timestep;
			signal=0.894154; #timestep;
			signal=0.892258; #timestep;
			signal=0.890349; #timestep;
			signal=0.888424; #timestep;
			signal=0.886485; #timestep;
			signal=0.884531; #timestep;
			signal=0.882563; #timestep;
			signal=0.88058; #timestep;
			signal=0.878583; #timestep;
			signal=0.876572; #timestep;
			signal=0.874546; #timestep;
			signal=0.872507; #timestep;
			signal=0.870453; #timestep;
			signal=0.868386; #timestep;
			signal=0.866305; #timestep;
			signal=0.864209; #timestep;
			signal=0.862101; #timestep;
			signal=0.859978; #timestep;
			signal=0.857842; #timestep;
			signal=0.855692; #timestep;
			signal=0.85353; #timestep;
			signal=0.851353; #timestep;
			signal=0.849164; #timestep;
			signal=0.846961; #timestep;
			signal=0.844746; #timestep;
			signal=0.842517; #timestep;
			signal=0.840275; #timestep;
			signal=0.838021; #timestep;
			signal=0.835754; #timestep;
			signal=0.833474; #timestep;
			signal=0.831182; #timestep;
			signal=0.828877; #timestep;
			signal=0.82656; #timestep;
			signal=0.824231; #timestep;
			signal=0.821889; #timestep;
			signal=0.819535; #timestep;
			signal=0.81717; #timestep;
			signal=0.814792; #timestep;
			signal=0.812402; #timestep;
			signal=0.810001; #timestep;
			signal=0.807588; #timestep;
			signal=0.805163; #timestep;
			signal=0.802727; #timestep;
			signal=0.80028; #timestep;
			signal=0.797821; #timestep;
			signal=0.795351; #timestep;
			signal=0.79287; #timestep;
			signal=0.790378; #timestep;
			signal=0.787875; #timestep;
			signal=0.785361; #timestep;
			signal=0.782836; #timestep;
			signal=0.780301; #timestep;
			signal=0.777755; #timestep;
			signal=0.775198; #timestep;
			signal=0.772632; #timestep;
			signal=0.770055; #timestep;
			signal=0.767468; #timestep;
			signal=0.76487; #timestep;
			signal=0.762263; #timestep;
			signal=0.759646; #timestep;
			signal=0.757019; #timestep;
			signal=0.754383; #timestep;
			signal=0.751737; #timestep;
			signal=0.749081; #timestep;
			signal=0.746416; #timestep;
			signal=0.743742; #timestep;
			signal=0.741059; #timestep;
			signal=0.738366; #timestep;
			signal=0.735665; #timestep;
			signal=0.732955; #timestep;
			signal=0.730236; #timestep;
			signal=0.727508; #timestep;
			signal=0.724771; #timestep;
			signal=0.722027; #timestep;
			signal=0.719274; #timestep;
			signal=0.716512; #timestep;
			signal=0.713743; #timestep;
			signal=0.710965; #timestep;
			signal=0.70818; #timestep;
			signal=0.705386; #timestep;
			signal=0.702585; #timestep;
			signal=0.699776; #timestep;
			signal=0.69696; #timestep;
			signal=0.694136; #timestep;
			signal=0.691305; #timestep;
			signal=0.688467; #timestep;
			signal=0.685622; #timestep;
			signal=0.68277; #timestep;
			signal=0.679911; #timestep;
			signal=0.677045; #timestep;
			signal=0.674172; #timestep;
			signal=0.671293; #timestep;
			signal=0.668407; #timestep;
			signal=0.665515; #timestep;
			signal=0.662617; #timestep;
			signal=0.659713; #timestep;
			signal=0.656803; #timestep;
			signal=0.653886; #timestep;
			signal=0.650964; #timestep;
			signal=0.648037; #timestep;
			signal=0.645103; #timestep;
			signal=0.642165; #timestep;
			signal=0.639221; #timestep;
			signal=0.636271; #timestep;
			signal=0.633317; #timestep;
			signal=0.630357; #timestep;
			signal=0.627393; #timestep;
			signal=0.624424; #timestep;
			signal=0.62145; #timestep;
			signal=0.618471; #timestep;
			signal=0.615489; #timestep;
			signal=0.612501; #timestep;
			signal=0.60951; #timestep;
			signal=0.606514; #timestep;
			signal=0.603515; #timestep;
			signal=0.600511; #timestep;
			signal=0.597504; #timestep;
			signal=0.594493; #timestep;
			signal=0.591478; #timestep;
			signal=0.58846; #timestep;
			signal=0.585439; #timestep;
			signal=0.582415; #timestep;
			signal=0.579387; #timestep;
			signal=0.576356; #timestep;
			signal=0.573323; #timestep;
			signal=0.570287; #timestep;
			signal=0.567248; #timestep;
			signal=0.564206; #timestep;
			signal=0.561162; #timestep;
			signal=0.558116; #timestep;
			signal=0.555068; #timestep;
			signal=0.552018; #timestep;
			signal=0.548965; #timestep;
			signal=0.545911; #timestep;
			signal=0.542855; #timestep;
			signal=0.539798; #timestep;
			signal=0.536739; #timestep;
			signal=0.533678; #timestep;
			signal=0.530616; #timestep;
			signal=0.527554; #timestep;
			signal=0.52449; #timestep;
			signal=0.521425; #timestep;
			signal=0.518359; #timestep;
			signal=0.515293; #timestep;
			signal=0.512226; #timestep;
			signal=0.509159; #timestep;
			signal=0.506091; #timestep;
			signal=0.503023; #timestep;
			signal=0.499955; #timestep;
			signal=0.496887; #timestep;
			signal=0.493819; #timestep;
			signal=0.490751; #timestep;
			signal=0.487684; #timestep;
			signal=0.484617; #timestep;
			signal=0.481551; #timestep;
			signal=0.478485; #timestep;
			signal=0.475421; #timestep;
			signal=0.472357; #timestep;
			signal=0.469294; #timestep;
			signal=0.466232; #timestep;
			signal=0.463172; #timestep;
			signal=0.460113; #timestep;
			signal=0.457055; #timestep;
			signal=0.453999; #timestep;
			signal=0.450945; #timestep;
			signal=0.447893; #timestep;
			signal=0.444843; #timestep;
			signal=0.441794; #timestep;
			signal=0.438748; #timestep;
			signal=0.435705; #timestep;
			signal=0.432663; #timestep;
			signal=0.429624; #timestep;
			signal=0.426588; #timestep;
			signal=0.423555; #timestep;
			signal=0.420524; #timestep;
			signal=0.417497; #timestep;
			signal=0.414472; #timestep;
			signal=0.411451; #timestep;
			signal=0.408433; #timestep;
			signal=0.405419; #timestep;
			signal=0.402408; #timestep;
			signal=0.399401; #timestep;
			signal=0.396397; #timestep;
			signal=0.393398; #timestep;
			signal=0.390402; #timestep;
			signal=0.387411; #timestep;
			signal=0.384424; #timestep;
			signal=0.381441; #timestep;
			signal=0.378463; #timestep;
			signal=0.375489; #timestep;
			signal=0.37252; #timestep;
			signal=0.369556; #timestep;
			signal=0.366597; #timestep;
			signal=0.363642; #timestep;
			signal=0.360693; #timestep;
			signal=0.357749; #timestep;
			signal=0.354811; #timestep;
			signal=0.351878; #timestep;
			signal=0.34895; #timestep;
			signal=0.346028; #timestep;
			signal=0.343112; #timestep;
			signal=0.340202; #timestep;
			signal=0.337298; #timestep;
			signal=0.3344; #timestep;
			signal=0.331508; #timestep;
			signal=0.328623; #timestep;
			signal=0.325744; #timestep;
			signal=0.322871; #timestep;
			signal=0.320006; #timestep;
			signal=0.317147; #timestep;
			signal=0.314295; #timestep;
			signal=0.31145; #timestep;
			signal=0.308612; #timestep;
			signal=0.305781; #timestep;
			signal=0.302957; #timestep;
			signal=0.300141; #timestep;
			signal=0.297333; #timestep;
			signal=0.294532; #timestep;
			signal=0.291739; #timestep;
			signal=0.288953; #timestep;
			signal=0.286176; #timestep;
			signal=0.283407; #timestep;
			signal=0.280646; #timestep;
			signal=0.277893; #timestep;
			signal=0.275148; #timestep;
			signal=0.272412; #timestep;
			signal=0.269685; #timestep;
			signal=0.266966; #timestep;
			signal=0.264256; #timestep;
			signal=0.261555; #timestep;
			signal=0.258862; #timestep;
			signal=0.256179; #timestep;
			signal=0.253505; #timestep;
			signal=0.250841; #timestep;
			signal=0.248185; #timestep;
			signal=0.24554; #timestep;
			signal=0.242903; #timestep;
			signal=0.240277; #timestep;
			signal=0.23766; #timestep;
			signal=0.235053; #timestep;
			signal=0.232456; #timestep;
			signal=0.22987; #timestep;
			signal=0.227293; #timestep;
			signal=0.224727; #timestep;
			signal=0.222171; #timestep;
			signal=0.219625; #timestep;
			signal=0.21709; #timestep;
			signal=0.214566; #timestep;
			signal=0.212052; #timestep;
			signal=0.209549; #timestep;
			signal=0.207057; #timestep;
			signal=0.204577; #timestep;
			signal=0.202107; #timestep;
			signal=0.199648; #timestep;
			signal=0.197201; #timestep;
			signal=0.194766; #timestep;
			signal=0.192341; #timestep;
			signal=0.189929; #timestep;
			signal=0.187528; #timestep;
			signal=0.185138; #timestep;
			signal=0.182761; #timestep;
			signal=0.180396; #timestep;
			signal=0.178042; #timestep;
			signal=0.175701; #timestep;
			signal=0.173372; #timestep;
			signal=0.171055; #timestep;
			signal=0.168751; #timestep;
			signal=0.166459; #timestep;
			signal=0.164179; #timestep;
			signal=0.161913; #timestep;
			signal=0.159659; #timestep;
			signal=0.157418; #timestep;
			signal=0.155189; #timestep;
			signal=0.152974; #timestep;
			signal=0.150772; #timestep;
			signal=0.148583; #timestep;
			signal=0.146407; #timestep;
			signal=0.144244; #timestep;
			signal=0.142095; #timestep;
			signal=0.13996; #timestep;
			signal=0.137837; #timestep;
			signal=0.135729; #timestep;
			signal=0.133634; #timestep;
			signal=0.131553; #timestep;
			signal=0.129486; #timestep;
			signal=0.127433; #timestep;
			signal=0.125394; #timestep;
			signal=0.123369; #timestep;
			signal=0.121358; #timestep;
			signal=0.119362; #timestep;
			signal=0.117379; #timestep;
			signal=0.115412; #timestep;
			signal=0.113458; #timestep;
			signal=0.111519; #timestep;
			signal=0.109595; #timestep;
			signal=0.107686; #timestep;
			signal=0.105791; #timestep;
			signal=0.103911; #timestep;
			signal=0.102046; #timestep;
			signal=0.100196; #timestep;
			signal=0.0983615; #timestep;
			signal=0.0965417; #timestep;
			signal=0.0947372; #timestep;
			signal=0.0929478; #timestep;
			signal=0.0911738; #timestep;
			signal=0.0894152; #timestep;
			signal=0.0876721; #timestep;
			signal=0.0859445; #timestep;
			signal=0.0842324; #timestep;
			signal=0.0825361; #timestep;
			signal=0.0808554; #timestep;
			signal=0.0791905; #timestep;
			signal=0.0775415; #timestep;
			signal=0.0759084; #timestep;
			signal=0.0742912; #timestep;
			signal=0.0726901; #timestep;
			signal=0.071105; #timestep;
			signal=0.0695361; #timestep;
			signal=0.0679834; #timestep;
			signal=0.066447; #timestep;
			signal=0.0649269; #timestep;
			signal=0.0634232; #timestep;
			signal=0.0619359; #timestep;
			signal=0.0604651; #timestep;
			signal=0.0590109; #timestep;
			signal=0.0575733; #timestep;
			signal=0.0561523; #timestep;
			signal=0.054748; #timestep;
			signal=0.0533605; #timestep;
			signal=0.0519899; #timestep;
			signal=0.0506361; #timestep;
			signal=0.0492992; #timestep;
			signal=0.0479792; #timestep;
			signal=0.0466763; #timestep;
			signal=0.0453905; #timestep;
			signal=0.0441218; #timestep;
			signal=0.0428702; #timestep;
			signal=0.0416359; #timestep;
			signal=0.0404188; #timestep;
			signal=0.039219; #timestep;
			signal=0.0380366; #timestep;
			signal=0.0368716; #timestep;
			signal=0.035724; #timestep;
			signal=0.0345938; #timestep;
			signal=0.0334812; #timestep;
			signal=0.0323862; #timestep;
			signal=0.0313088; #timestep;
			signal=0.030249; #timestep;
			signal=0.0292069; #timestep;
			signal=0.0281826; #timestep;
			signal=0.027176; #timestep;
			signal=0.0261872; #timestep;
			signal=0.0252162; #timestep;
			signal=0.0242631; #timestep;
			signal=0.023328; #timestep;
			signal=0.0224107; #timestep;
			signal=0.0215115; #timestep;
			signal=0.0206303; #timestep;
			signal=0.0197671; #timestep;
			signal=0.018922; #timestep;
			signal=0.018095; #timestep;
			signal=0.0172862; #timestep;
			signal=0.0164955; #timestep;
			signal=0.0157231; #timestep;
			signal=0.0149689; #timestep;
			signal=0.0142329; #timestep;
			signal=0.0135152; #timestep;
			signal=0.0128159; #timestep;
			signal=0.0121349; #timestep;
			signal=0.0114722; #timestep;
			signal=0.010828; #timestep;
			signal=0.0102021; #timestep;
			signal=0.00959476; #timestep;
			signal=0.00900584; #timestep;
			signal=0.00843541; #timestep;
			signal=0.00788348; #timestep;
			signal=0.00735008; #timestep;
			signal=0.00683523; #timestep;
			signal=0.00633895; #timestep;
			signal=0.00586126; #timestep;
			signal=0.00540217; #timestep;
			signal=0.0049617; #timestep;
			signal=0.00453988; #timestep;
			signal=0.0041367; #timestep;
			signal=0.0037522; #timestep;
			signal=0.00338638; #timestep;
			signal=0.00303926; #timestep;
			signal=0.00271086; #timestep;
			signal=0.00240117; #timestep;
			signal=0.00211022; #timestep;
			signal=0.00183802; #timestep;
			signal=0.00158458; #timestep;
			signal=0.0013499; #timestep;
			signal=0.00113399; #timestep;
			signal=0.000936869; #timestep;
			signal=0.000758538; #timestep;
			signal=0.000599004; #timestep;
			signal=0.000458273; #timestep;
			signal=0.000336351; #timestep;
			signal=0.000233242; #timestep;
			signal=0.00014895; #timestep;
			signal=8.34779e-005; #timestep;
			signal=3.68287e-005; #timestep;
			signal=9.00388e-006; #timestep;
			signal=4.54256e-009; #timestep;
			signal=9.831e-006; #timestep;
			signal=3.84829e-005; #timestep;
			signal=8.59591e-005; #timestep;
			signal=0.000152258; #timestep;
			signal=0.000237377; #timestep;
			signal=0.000341312; #timestep;
			signal=0.000464061; #timestep;
			signal=0.000605618; #timestep;
			signal=0.000765978; #timestep;
			signal=0.000945135; #timestep;
			signal=0.00114308; #timestep;
			signal=0.00135981; #timestep;
			signal=0.00159532; #timestep;
			signal=0.00184959; #timestep;
			signal=0.00212261; #timestep;
			signal=0.00241439; #timestep;
			signal=0.00272489; #timestep;
			signal=0.00305412; #timestep;
			signal=0.00340206; #timestep;
			signal=0.0037687; #timestep;
			signal=0.00415403; #timestep;
			signal=0.00455802; #timestep;
			signal=0.00498066; #timestep;
			signal=0.00542195; #timestep;
			signal=0.00588185; #timestep;
			signal=0.00636036; #timestep;
			signal=0.00685746; #timestep;
			signal=0.00737313; #timestep;
			signal=0.00790734; #timestep;
			signal=0.00846008; #timestep;
			signal=0.00903133; #timestep;
			signal=0.00962106; #timestep;
			signal=0.0102293; #timestep;
			signal=0.0108559; #timestep;
			signal=0.011501; #timestep;
			signal=0.0121644; #timestep;
			signal=0.0128462; #timestep;
			signal=0.0135464; #timestep;
			signal=0.0142648; #timestep;
			signal=0.0150016; #timestep;
			signal=0.0157566; #timestep;
			signal=0.0165299; #timestep;
			signal=0.0173213; #timestep;
			signal=0.018131; #timestep;
			signal=0.0189588; #timestep;
			signal=0.0198046; #timestep;
			signal=0.0206686; #timestep;
			signal=0.0215506; #timestep;
			signal=0.0224507; #timestep;
			signal=0.0233687; #timestep;
			signal=0.0243046; #timestep;
			signal=0.0252585; #timestep;
			signal=0.0262302; #timestep;
			signal=0.0272198; #timestep;
			signal=0.0282272; #timestep;
			signal=0.0292523; #timestep;
			signal=0.0302952; #timestep;
			signal=0.0313558; #timestep;
			signal=0.032434; #timestep;
			signal=0.0335298; #timestep;
			signal=0.0346431; #timestep;
			signal=0.035774; #timestep;
			signal=0.0369224; #timestep;
			signal=0.0380882; #timestep;
			signal=0.0392714; #timestep;
			signal=0.0404719; #timestep;
			signal=0.0416898; #timestep;
			signal=0.0429249; #timestep;
			signal=0.0441772; #timestep;
			signal=0.0454466; #timestep;
			signal=0.0467332; #timestep;
			signal=0.0480369; #timestep;
			signal=0.0493575; #timestep;
			signal=0.0506952; #timestep;
			signal=0.0520497; #timestep;
			signal=0.0534212; #timestep;
			signal=0.0548094; #timestep;
			signal=0.0562144; #timestep;
			signal=0.0576361; #timestep;
			signal=0.0590745; #timestep;
			signal=0.0605294; #timestep;
			signal=0.0620009; #timestep;
			signal=0.0634889; #timestep;
			signal=0.0649934; #timestep;
			signal=0.0665142; #timestep;
			signal=0.0680513; #timestep;
			signal=0.0696047; #timestep;
			signal=0.0711743; #timestep;
			signal=0.0727601; #timestep;
			signal=0.0743619; #timestep;
			signal=0.0759798; #timestep;
			signal=0.0776136; #timestep;
			signal=0.0792633; #timestep;
			signal=0.0809289; #timestep;
			signal=0.0826103; #timestep;
			signal=0.0843073; #timestep;
			signal=0.08602; #timestep;
			signal=0.0877483; #timestep;
			signal=0.0894922; #timestep;
			signal=0.0912515; #timestep;
			signal=0.0930261; #timestep;
			signal=0.0948161; #timestep;
			signal=0.0966214; #timestep;
			signal=0.0984418; #timestep;
			signal=0.100277; #timestep;
			signal=0.102128; #timestep;
			signal=0.103994; #timestep;
			signal=0.105874; #timestep;
			signal=0.107769; #timestep;
			signal=0.10968; #timestep;
			signal=0.111604; #timestep;
			signal=0.113544; #timestep;
			signal=0.115498; #timestep;
			signal=0.117466; #timestep;
			signal=0.119449; #timestep;
			signal=0.121446; #timestep;
			signal=0.123458; #timestep;
			signal=0.125483; #timestep;
			signal=0.127523; #timestep;
			signal=0.129577; #timestep;
			signal=0.131644; #timestep;
			signal=0.133726; #timestep;
			signal=0.135821; #timestep;
			signal=0.13793; #timestep;
			signal=0.140053; #timestep;
			signal=0.142189; #timestep;
			signal=0.144339; #timestep;
			signal=0.146502; #timestep;
			signal=0.148679; #timestep;
			signal=0.150868; #timestep;
			signal=0.153071; #timestep;
			signal=0.155287; #timestep;
			signal=0.157516; #timestep;
			signal=0.159758; #timestep;
			signal=0.162012; #timestep;
			signal=0.164279; #timestep;
			signal=0.166559; #timestep;
			signal=0.168852; #timestep;
			signal=0.171157; #timestep;
			signal=0.173474; #timestep;
			signal=0.175804; #timestep;
			signal=0.178145; #timestep;
			signal=0.180499; #timestep;
			signal=0.182865; #timestep;
			signal=0.185243; #timestep;
			signal=0.187633; #timestep;
			signal=0.190034; #timestep;
			signal=0.192448; #timestep;
			signal=0.194872; #timestep;
			signal=0.197309; #timestep;
			signal=0.199756; #timestep;
			signal=0.202215; #timestep;
			signal=0.204685; #timestep;
			signal=0.207167; #timestep;
			signal=0.209659; #timestep;
			signal=0.212162; #timestep;
			signal=0.214676; #timestep;
			signal=0.217201; #timestep;
			signal=0.219737; #timestep;
			signal=0.222283; #timestep;
			signal=0.224839; #timestep;
			signal=0.227406; #timestep;
			signal=0.229983; #timestep;
			signal=0.23257; #timestep;
			signal=0.235168; #timestep;
			signal=0.237775; #timestep;
			signal=0.240392; #timestep;
			signal=0.243019; #timestep;
			signal=0.245656; #timestep;
			signal=0.248302; #timestep;
			signal=0.250958; #timestep;
			signal=0.253623; #timestep;
			signal=0.256297; #timestep;
			signal=0.258981; #timestep;
			signal=0.261673; #timestep;
			signal=0.264375; #timestep;
			signal=0.267085; #timestep;
			signal=0.269804; #timestep;
			signal=0.272532; #timestep;
			signal=0.275269; #timestep;
			signal=0.278014; #timestep;
			signal=0.280767; #timestep;
			signal=0.283528; #timestep;
			signal=0.286298; #timestep;
			signal=0.289076; #timestep;
			signal=0.291861; #timestep;
			signal=0.294655; #timestep;
			signal=0.297456; #timestep;
			signal=0.300265; #timestep;
			signal=0.303081; #timestep;
			signal=0.305905; #timestep;
			signal=0.308736; #timestep;
			signal=0.311574; #timestep;
			signal=0.31442; #timestep;
			signal=0.317272; #timestep;
			signal=0.320131; #timestep;
			signal=0.322997; #timestep;
			signal=0.32587; #timestep;
			signal=0.328749; #timestep;
			signal=0.331635; #timestep;
			signal=0.334527; #timestep;
			signal=0.337425; #timestep;
			signal=0.34033; #timestep;
			signal=0.34324; #timestep;
			signal=0.346156; #timestep;
			signal=0.349079; #timestep;
			signal=0.352006; #timestep;
			signal=0.35494; #timestep;
			signal=0.357878; #timestep;
			signal=0.360823; #timestep;
			signal=0.363772; #timestep;
			signal=0.366727; #timestep;
			signal=0.369686; #timestep;
			signal=0.372651; #timestep;
			signal=0.37562; #timestep;
			signal=0.378594; #timestep;
			signal=0.381572; #timestep;
			signal=0.384555; #timestep;
			signal=0.387542; #timestep;
			signal=0.390534; #timestep;
			signal=0.39353; #timestep;
			signal=0.396529; #timestep;
			signal=0.399533; #timestep;
			signal=0.40254; #timestep;
			signal=0.405551; #timestep;
			signal=0.408566; #timestep;
			signal=0.411584; #timestep;
			signal=0.414605; #timestep;
			signal=0.41763; #timestep;
			signal=0.420657; #timestep;
			signal=0.423688; #timestep;
			signal=0.426722; #timestep;
			signal=0.429758; #timestep;
			signal=0.432797; #timestep;
			signal=0.435838; #timestep;
			signal=0.438882; #timestep;
			signal=0.441928; #timestep;
			signal=0.444977; #timestep;
			signal=0.448027; #timestep;
			signal=0.451079; #timestep;
			signal=0.454134; #timestep;
			signal=0.45719; #timestep;
			signal=0.460247; #timestep;
			signal=0.463306; #timestep;
			signal=0.466367; #timestep;
			signal=0.469428; #timestep;
			signal=0.472491; #timestep;
			signal=0.475555; #timestep;
			signal=0.47862; #timestep;
			signal=0.481686; #timestep;
			signal=0.484752; #timestep;
			signal=0.487819; #timestep;
			signal=0.490886; #timestep;
			signal=0.493954; #timestep;
			signal=0.497022; #timestep;
		end 
endmodule