// one module to rule them all...

module topModule (
    input logic [1:0] ps2keyBoard,
    input logic [7:0] buttonBoard,
    input logic clk,
    output logic [6:0] segments
    );

    // its 3 am... im going to bed

endmodule